module mux_256x32b_to_1x32b (out, in, select);

  output [31:0] out;
  input [32767:0] in;
  input [9:0] select; //read address now 10 bits long for 1024 locations

  reg [31:0] out;

  always @ (in or select) begin
    casex(select)
// %%start_veriperl
// my $i;
// my $low_index;
// my $high_index;
// for($i=0; $i<1024; $i=$i+1)
// {
//   $low_index = 32*$i;
//   $high_index = 32*$i+31;
//   print "      10'd$i : out <= in [$high_index:$low_index];\n";
// }
// %%stop_veriperl
      10'd0 : out <= in [31:0];
      10'd1 : out <= in [63:32];
      10'd2 : out <= in [95:64];
      10'd3 : out <= in [127:96];
      10'd4 : out <= in [159:128];
      10'd5 : out <= in [191:160];
      10'd6 : out <= in [223:192];
      10'd7 : out <= in [255:224];
      10'd8 : out <= in [287:256];
      10'd9 : out <= in [319:288];
      10'd10 : out <= in [351:320];
      10'd11 : out <= in [383:352];
      10'd12 : out <= in [415:384];
      10'd13 : out <= in [447:416];
      10'd14 : out <= in [479:448];
      10'd15 : out <= in [511:480];
      10'd16 : out <= in [543:512];
      10'd17 : out <= in [575:544];
      10'd18 : out <= in [607:576];
      10'd19 : out <= in [639:608];
      10'd20 : out <= in [671:640];
      10'd21 : out <= in [703:672];
      10'd22 : out <= in [735:704];
      10'd23 : out <= in [767:736];
      10'd24 : out <= in [799:768];
      10'd25 : out <= in [831:800];
      10'd26 : out <= in [863:832];
      10'd27 : out <= in [895:864];
      10'd28 : out <= in [927:896];
      10'd29 : out <= in [959:928];
      10'd30 : out <= in [991:960];
      10'd31 : out <= in [1023:992];
      10'd32 : out <= in [1055:1024];
      10'd33 : out <= in [1087:1056];
      10'd34 : out <= in [1119:1088];
      10'd35 : out <= in [1151:1120];
      10'd36 : out <= in [1183:1152];
      10'd37 : out <= in [1215:1184];
      10'd38 : out <= in [1247:1216];
      10'd39 : out <= in [1279:1248];
      10'd40 : out <= in [1311:1280];
      10'd41 : out <= in [1343:1312];
      10'd42 : out <= in [1375:1344];
      10'd43 : out <= in [1407:1376];
      10'd44 : out <= in [1439:1408];
      10'd45 : out <= in [1471:1440];
      10'd46 : out <= in [1503:1472];
      10'd47 : out <= in [1535:1504];
      10'd48 : out <= in [1567:1536];
      10'd49 : out <= in [1599:1568];
      10'd50 : out <= in [1631:1600];
      10'd51 : out <= in [1663:1632];
      10'd52 : out <= in [1695:1664];
      10'd53 : out <= in [1727:1696];
      10'd54 : out <= in [1759:1728];
      10'd55 : out <= in [1791:1760];
      10'd56 : out <= in [1823:1792];
      10'd57 : out <= in [1855:1824];
      10'd58 : out <= in [1887:1856];
      10'd59 : out <= in [1919:1888];
      10'd60 : out <= in [1951:1920];
      10'd61 : out <= in [1983:1952];
      10'd62 : out <= in [2015:1984];
      10'd63 : out <= in [2047:2016];
      10'd64 : out <= in [2079:2048];
      10'd65 : out <= in [2111:2080];
      10'd66 : out <= in [2143:2112];
      10'd67 : out <= in [2175:2144];
      10'd68 : out <= in [2207:2176];
      10'd69 : out <= in [2239:2208];
      10'd70 : out <= in [2271:2240];
      10'd71 : out <= in [2303:2272];
      10'd72 : out <= in [2335:2304];
      10'd73 : out <= in [2367:2336];
      10'd74 : out <= in [2399:2368];
      10'd75 : out <= in [2431:2400];
      10'd76 : out <= in [2463:2432];
      10'd77 : out <= in [2495:2464];
      10'd78 : out <= in [2527:2496];
      10'd79 : out <= in [2559:2528];
      10'd80 : out <= in [2591:2560];
      10'd81 : out <= in [2623:2592];
      10'd82 : out <= in [2655:2624];
      10'd83 : out <= in [2687:2656];
      10'd84 : out <= in [2719:2688];
      10'd85 : out <= in [2751:2720];
      10'd86 : out <= in [2783:2752];
      10'd87 : out <= in [2815:2784];
      10'd88 : out <= in [2847:2816];
      10'd89 : out <= in [2879:2848];
      10'd90 : out <= in [2911:2880];
      10'd91 : out <= in [2943:2912];
      10'd92 : out <= in [2975:2944];
      10'd93 : out <= in [3007:2976];
      10'd94 : out <= in [3039:3008];
      10'd95 : out <= in [3071:3040];
      10'd96 : out <= in [3103:3072];
      10'd97 : out <= in [3135:3104];
      10'd98 : out <= in [3167:3136];
      10'd99 : out <= in [3199:3168];
      10'd100 : out <= in [3231:3200];
      10'd101 : out <= in [3263:3232];
      10'd102 : out <= in [3295:3264];
      10'd103 : out <= in [3327:3296];
      10'd104 : out <= in [3359:3328];
      10'd105 : out <= in [3391:3360];
      10'd106 : out <= in [3423:3392];
      10'd107 : out <= in [3455:3424];
      10'd108 : out <= in [3487:3456];
      10'd109 : out <= in [3519:3488];
      10'd110 : out <= in [3551:3520];
      10'd111 : out <= in [3583:3552];
      10'd112 : out <= in [3615:3584];
      10'd113 : out <= in [3647:3616];
      10'd114 : out <= in [3679:3648];
      10'd115 : out <= in [3711:3680];
      10'd116 : out <= in [3743:3712];
      10'd117 : out <= in [3775:3744];
      10'd118 : out <= in [3807:3776];
      10'd119 : out <= in [3839:3808];
      10'd120 : out <= in [3871:3840];
      10'd121 : out <= in [3903:3872];
      10'd122 : out <= in [3935:3904];
      10'd123 : out <= in [3967:3936];
      10'd124 : out <= in [3999:3968];
      10'd125 : out <= in [4031:4000];
      10'd126 : out <= in [4063:4032];
      10'd127 : out <= in [4095:4064];
      10'd128 : out <= in [4127:4096];
      10'd129 : out <= in [4159:4128];
      10'd130 : out <= in [4191:4160];
      10'd131 : out <= in [4223:4192];
      10'd132 : out <= in [4255:4224];
      10'd133 : out <= in [4287:4256];
      10'd134 : out <= in [4319:4288];
      10'd135 : out <= in [4351:4320];
      10'd136 : out <= in [4383:4352];
      10'd137 : out <= in [4415:4384];
      10'd138 : out <= in [4447:4416];
      10'd139 : out <= in [4479:4448];
      10'd140 : out <= in [4511:4480];
      10'd141 : out <= in [4543:4512];
      10'd142 : out <= in [4575:4544];
      10'd143 : out <= in [4607:4576];
      10'd144 : out <= in [4639:4608];
      10'd145 : out <= in [4671:4640];
      10'd146 : out <= in [4703:4672];
      10'd147 : out <= in [4735:4704];
      10'd148 : out <= in [4767:4736];
      10'd149 : out <= in [4799:4768];
      10'd150 : out <= in [4831:4800];
      10'd151 : out <= in [4863:4832];
      10'd152 : out <= in [4895:4864];
      10'd153 : out <= in [4927:4896];
      10'd154 : out <= in [4959:4928];
      10'd155 : out <= in [4991:4960];
      10'd156 : out <= in [5023:4992];
      10'd157 : out <= in [5055:5024];
      10'd158 : out <= in [5087:5056];
      10'd159 : out <= in [5119:5088];
      10'd160 : out <= in [5151:5120];
      10'd161 : out <= in [5183:5152];
      10'd162 : out <= in [5215:5184];
      10'd163 : out <= in [5247:5216];
      10'd164 : out <= in [5279:5248];
      10'd165 : out <= in [5311:5280];
      10'd166 : out <= in [5343:5312];
      10'd167 : out <= in [5375:5344];
      10'd168 : out <= in [5407:5376];
      10'd169 : out <= in [5439:5408];
      10'd170 : out <= in [5471:5440];
      10'd171 : out <= in [5503:5472];
      10'd172 : out <= in [5535:5504];
      10'd173 : out <= in [5567:5536];
      10'd174 : out <= in [5599:5568];
      10'd175 : out <= in [5631:5600];
      10'd176 : out <= in [5663:5632];
      10'd177 : out <= in [5695:5664];
      10'd178 : out <= in [5727:5696];
      10'd179 : out <= in [5759:5728];
      10'd180 : out <= in [5791:5760];
      10'd181 : out <= in [5823:5792];
      10'd182 : out <= in [5855:5824];
      10'd183 : out <= in [5887:5856];
      10'd184 : out <= in [5919:5888];
      10'd185 : out <= in [5951:5920];
      10'd186 : out <= in [5983:5952];
      10'd187 : out <= in [6015:5984];
      10'd188 : out <= in [6047:6016];
      10'd189 : out <= in [6079:6048];
      10'd190 : out <= in [6111:6080];
      10'd191 : out <= in [6143:6112];
      10'd192 : out <= in [6175:6144];
      10'd193 : out <= in [6207:6176];
      10'd194 : out <= in [6239:6208];
      10'd195 : out <= in [6271:6240];
      10'd196 : out <= in [6303:6272];
      10'd197 : out <= in [6335:6304];
      10'd198 : out <= in [6367:6336];
      10'd199 : out <= in [6399:6368];
      10'd200 : out <= in [6431:6400];
      10'd201 : out <= in [6463:6432];
      10'd202 : out <= in [6495:6464];
      10'd203 : out <= in [6527:6496];
      10'd204 : out <= in [6559:6528];
      10'd205 : out <= in [6591:6560];
      10'd206 : out <= in [6623:6592];
      10'd207 : out <= in [6655:6624];
      10'd208 : out <= in [6687:6656];
      10'd209 : out <= in [6719:6688];
      10'd210 : out <= in [6751:6720];
      10'd211 : out <= in [6783:6752];
      10'd212 : out <= in [6815:6784];
      10'd213 : out <= in [6847:6816];
      10'd214 : out <= in [6879:6848];
      10'd215 : out <= in [6911:6880];
      10'd216 : out <= in [6943:6912];
      10'd217 : out <= in [6975:6944];
      10'd218 : out <= in [7007:6976];
      10'd219 : out <= in [7039:7008];
      10'd220 : out <= in [7071:7040];
      10'd221 : out <= in [7103:7072];
      10'd222 : out <= in [7135:7104];
      10'd223 : out <= in [7167:7136];
      10'd224 : out <= in [7199:7168];
      10'd225 : out <= in [7231:7200];
      10'd226 : out <= in [7263:7232];
      10'd227 : out <= in [7295:7264];
      10'd228 : out <= in [7327:7296];
      10'd229 : out <= in [7359:7328];
      10'd230 : out <= in [7391:7360];
      10'd231 : out <= in [7423:7392];
      10'd232 : out <= in [7455:7424];
      10'd233 : out <= in [7487:7456];
      10'd234 : out <= in [7519:7488];
      10'd235 : out <= in [7551:7520];
      10'd236 : out <= in [7583:7552];
      10'd237 : out <= in [7615:7584];
      10'd238 : out <= in [7647:7616];
      10'd239 : out <= in [7679:7648];
      10'd240 : out <= in [7711:7680];
      10'd241 : out <= in [7743:7712];
      10'd242 : out <= in [7775:7744];
      10'd243 : out <= in [7807:7776];
      10'd244 : out <= in [7839:7808];
      10'd245 : out <= in [7871:7840];
      10'd246 : out <= in [7903:7872];
      10'd247 : out <= in [7935:7904];
      10'd248 : out <= in [7967:7936];
      10'd249 : out <= in [7999:7968];
      10'd250 : out <= in [8031:8000];
      10'd251 : out <= in [8063:8032];
      10'd252 : out <= in [8095:8064];
      10'd253 : out <= in [8127:8096];
      10'd254 : out <= in [8159:8128];
      10'd255 : out <= in [8191:8160];
      10'd256 : out <= in [8223:8192];
      10'd257 : out <= in [8255:8224];
      10'd258 : out <= in [8287:8256];
      10'd259 : out <= in [8319:8288];
      10'd260 : out <= in [8351:8320];
      10'd261 : out <= in [8383:8352];
      10'd262 : out <= in [8415:8384];
      10'd263 : out <= in [8447:8416];
      10'd264 : out <= in [8479:8448];
      10'd265 : out <= in [8511:8480];
      10'd266 : out <= in [8543:8512];
      10'd267 : out <= in [8575:8544];
      10'd268 : out <= in [8607:8576];
      10'd269 : out <= in [8639:8608];
      10'd270 : out <= in [8671:8640];
      10'd271 : out <= in [8703:8672];
      10'd272 : out <= in [8735:8704];
      10'd273 : out <= in [8767:8736];
      10'd274 : out <= in [8799:8768];
      10'd275 : out <= in [8831:8800];
      10'd276 : out <= in [8863:8832];
      10'd277 : out <= in [8895:8864];
      10'd278 : out <= in [8927:8896];
      10'd279 : out <= in [8959:8928];
      10'd280 : out <= in [8991:8960];
      10'd281 : out <= in [9023:8992];
      10'd282 : out <= in [9055:9024];
      10'd283 : out <= in [9087:9056];
      10'd284 : out <= in [9119:9088];
      10'd285 : out <= in [9151:9120];
      10'd286 : out <= in [9183:9152];
      10'd287 : out <= in [9215:9184];
      10'd288 : out <= in [9247:9216];
      10'd289 : out <= in [9279:9248];
      10'd290 : out <= in [9311:9280];
      10'd291 : out <= in [9343:9312];
      10'd292 : out <= in [9375:9344];
      10'd293 : out <= in [9407:9376];
      10'd294 : out <= in [9439:9408];
      10'd295 : out <= in [9471:9440];
      10'd296 : out <= in [9503:9472];
      10'd297 : out <= in [9535:9504];
      10'd298 : out <= in [9567:9536];
      10'd299 : out <= in [9599:9568];
      10'd300 : out <= in [9631:9600];
      10'd301 : out <= in [9663:9632];
      10'd302 : out <= in [9695:9664];
      10'd303 : out <= in [9727:9696];
      10'd304 : out <= in [9759:9728];
      10'd305 : out <= in [9791:9760];
      10'd306 : out <= in [9823:9792];
      10'd307 : out <= in [9855:9824];
      10'd308 : out <= in [9887:9856];
      10'd309 : out <= in [9919:9888];
      10'd310 : out <= in [9951:9920];
      10'd311 : out <= in [9983:9952];
      10'd312 : out <= in [10015:9984];
      10'd313 : out <= in [10047:10016];
      10'd314 : out <= in [10079:10048];
      10'd315 : out <= in [10111:10080];
      10'd316 : out <= in [10143:10112];
      10'd317 : out <= in [10175:10144];
      10'd318 : out <= in [10207:10176];
      10'd319 : out <= in [10239:10208];
      10'd320 : out <= in [10271:10240];
      10'd321 : out <= in [10303:10272];
      10'd322 : out <= in [10335:10304];
      10'd323 : out <= in [10367:10336];
      10'd324 : out <= in [10399:10368];
      10'd325 : out <= in [10431:10400];
      10'd326 : out <= in [10463:10432];
      10'd327 : out <= in [10495:10464];
      10'd328 : out <= in [10527:10496];
      10'd329 : out <= in [10559:10528];
      10'd330 : out <= in [10591:10560];
      10'd331 : out <= in [10623:10592];
      10'd332 : out <= in [10655:10624];
      10'd333 : out <= in [10687:10656];
      10'd334 : out <= in [10719:10688];
      10'd335 : out <= in [10751:10720];
      10'd336 : out <= in [10783:10752];
      10'd337 : out <= in [10815:10784];
      10'd338 : out <= in [10847:10816];
      10'd339 : out <= in [10879:10848];
      10'd340 : out <= in [10911:10880];
      10'd341 : out <= in [10943:10912];
      10'd342 : out <= in [10975:10944];
      10'd343 : out <= in [11007:10976];
      10'd344 : out <= in [11039:11008];
      10'd345 : out <= in [11071:11040];
      10'd346 : out <= in [11103:11072];
      10'd347 : out <= in [11135:11104];
      10'd348 : out <= in [11167:11136];
      10'd349 : out <= in [11199:11168];
      10'd350 : out <= in [11231:11200];
      10'd351 : out <= in [11263:11232];
      10'd352 : out <= in [11295:11264];
      10'd353 : out <= in [11327:11296];
      10'd354 : out <= in [11359:11328];
      10'd355 : out <= in [11391:11360];
      10'd356 : out <= in [11423:11392];
      10'd357 : out <= in [11455:11424];
      10'd358 : out <= in [11487:11456];
      10'd359 : out <= in [11519:11488];
      10'd360 : out <= in [11551:11520];
      10'd361 : out <= in [11583:11552];
      10'd362 : out <= in [11615:11584];
      10'd363 : out <= in [11647:11616];
      10'd364 : out <= in [11679:11648];
      10'd365 : out <= in [11711:11680];
      10'd366 : out <= in [11743:11712];
      10'd367 : out <= in [11775:11744];
      10'd368 : out <= in [11807:11776];
      10'd369 : out <= in [11839:11808];
      10'd370 : out <= in [11871:11840];
      10'd371 : out <= in [11903:11872];
      10'd372 : out <= in [11935:11904];
      10'd373 : out <= in [11967:11936];
      10'd374 : out <= in [11999:11968];
      10'd375 : out <= in [12031:12000];
      10'd376 : out <= in [12063:12032];
      10'd377 : out <= in [12095:12064];
      10'd378 : out <= in [12127:12096];
      10'd379 : out <= in [12159:12128];
      10'd380 : out <= in [12191:12160];
      10'd381 : out <= in [12223:12192];
      10'd382 : out <= in [12255:12224];
      10'd383 : out <= in [12287:12256];
      10'd384 : out <= in [12319:12288];
      10'd385 : out <= in [12351:12320];
      10'd386 : out <= in [12383:12352];
      10'd387 : out <= in [12415:12384];
      10'd388 : out <= in [12447:12416];
      10'd389 : out <= in [12479:12448];
      10'd390 : out <= in [12511:12480];
      10'd391 : out <= in [12543:12512];
      10'd392 : out <= in [12575:12544];
      10'd393 : out <= in [12607:12576];
      10'd394 : out <= in [12639:12608];
      10'd395 : out <= in [12671:12640];
      10'd396 : out <= in [12703:12672];
      10'd397 : out <= in [12735:12704];
      10'd398 : out <= in [12767:12736];
      10'd399 : out <= in [12799:12768];
      10'd400 : out <= in [12831:12800];
      10'd401 : out <= in [12863:12832];
      10'd402 : out <= in [12895:12864];
      10'd403 : out <= in [12927:12896];
      10'd404 : out <= in [12959:12928];
      10'd405 : out <= in [12991:12960];
      10'd406 : out <= in [13023:12992];
      10'd407 : out <= in [13055:13024];
      10'd408 : out <= in [13087:13056];
      10'd409 : out <= in [13119:13088];
      10'd410 : out <= in [13151:13120];
      10'd411 : out <= in [13183:13152];
      10'd412 : out <= in [13215:13184];
      10'd413 : out <= in [13247:13216];
      10'd414 : out <= in [13279:13248];
      10'd415 : out <= in [13311:13280];
      10'd416 : out <= in [13343:13312];
      10'd417 : out <= in [13375:13344];
      10'd418 : out <= in [13407:13376];
      10'd419 : out <= in [13439:13408];
      10'd420 : out <= in [13471:13440];
      10'd421 : out <= in [13503:13472];
      10'd422 : out <= in [13535:13504];
      10'd423 : out <= in [13567:13536];
      10'd424 : out <= in [13599:13568];
      10'd425 : out <= in [13631:13600];
      10'd426 : out <= in [13663:13632];
      10'd427 : out <= in [13695:13664];
      10'd428 : out <= in [13727:13696];
      10'd429 : out <= in [13759:13728];
      10'd430 : out <= in [13791:13760];
      10'd431 : out <= in [13823:13792];
      10'd432 : out <= in [13855:13824];
      10'd433 : out <= in [13887:13856];
      10'd434 : out <= in [13919:13888];
      10'd435 : out <= in [13951:13920];
      10'd436 : out <= in [13983:13952];
      10'd437 : out <= in [14015:13984];
      10'd438 : out <= in [14047:14016];
      10'd439 : out <= in [14079:14048];
      10'd440 : out <= in [14111:14080];
      10'd441 : out <= in [14143:14112];
      10'd442 : out <= in [14175:14144];
      10'd443 : out <= in [14207:14176];
      10'd444 : out <= in [14239:14208];
      10'd445 : out <= in [14271:14240];
      10'd446 : out <= in [14303:14272];
      10'd447 : out <= in [14335:14304];
      10'd448 : out <= in [14367:14336];
      10'd449 : out <= in [14399:14368];
      10'd450 : out <= in [14431:14400];
      10'd451 : out <= in [14463:14432];
      10'd452 : out <= in [14495:14464];
      10'd453 : out <= in [14527:14496];
      10'd454 : out <= in [14559:14528];
      10'd455 : out <= in [14591:14560];
      10'd456 : out <= in [14623:14592];
      10'd457 : out <= in [14655:14624];
      10'd458 : out <= in [14687:14656];
      10'd459 : out <= in [14719:14688];
      10'd460 : out <= in [14751:14720];
      10'd461 : out <= in [14783:14752];
      10'd462 : out <= in [14815:14784];
      10'd463 : out <= in [14847:14816];
      10'd464 : out <= in [14879:14848];
      10'd465 : out <= in [14911:14880];
      10'd466 : out <= in [14943:14912];
      10'd467 : out <= in [14975:14944];
      10'd468 : out <= in [15007:14976];
      10'd469 : out <= in [15039:15008];
      10'd470 : out <= in [15071:15040];
      10'd471 : out <= in [15103:15072];
      10'd472 : out <= in [15135:15104];
      10'd473 : out <= in [15167:15136];
      10'd474 : out <= in [15199:15168];
      10'd475 : out <= in [15231:15200];
      10'd476 : out <= in [15263:15232];
      10'd477 : out <= in [15295:15264];
      10'd478 : out <= in [15327:15296];
      10'd479 : out <= in [15359:15328];
      10'd480 : out <= in [15391:15360];
      10'd481 : out <= in [15423:15392];
      10'd482 : out <= in [15455:15424];
      10'd483 : out <= in [15487:15456];
      10'd484 : out <= in [15519:15488];
      10'd485 : out <= in [15551:15520];
      10'd486 : out <= in [15583:15552];
      10'd487 : out <= in [15615:15584];
      10'd488 : out <= in [15647:15616];
      10'd489 : out <= in [15679:15648];
      10'd490 : out <= in [15711:15680];
      10'd491 : out <= in [15743:15712];
      10'd492 : out <= in [15775:15744];
      10'd493 : out <= in [15807:15776];
      10'd494 : out <= in [15839:15808];
      10'd495 : out <= in [15871:15840];
      10'd496 : out <= in [15903:15872];
      10'd497 : out <= in [15935:15904];
      10'd498 : out <= in [15967:15936];
      10'd499 : out <= in [15999:15968];
      10'd500 : out <= in [16031:16000];
      10'd501 : out <= in [16063:16032];
      10'd502 : out <= in [16095:16064];
      10'd503 : out <= in [16127:16096];
      10'd504 : out <= in [16159:16128];
      10'd505 : out <= in [16191:16160];
      10'd506 : out <= in [16223:16192];
      10'd507 : out <= in [16255:16224];
      10'd508 : out <= in [16287:16256];
      10'd509 : out <= in [16319:16288];
      10'd510 : out <= in [16351:16320];
      10'd511 : out <= in [16383:16352];
      10'd512 : out <= in [16415:16384];
      10'd513 : out <= in [16447:16416];
      10'd514 : out <= in [16479:16448];
      10'd515 : out <= in [16511:16480];
      10'd516 : out <= in [16543:16512];
      10'd517 : out <= in [16575:16544];
      10'd518 : out <= in [16607:16576];
      10'd519 : out <= in [16639:16608];
      10'd520 : out <= in [16671:16640];
      10'd521 : out <= in [16703:16672];
      10'd522 : out <= in [16735:16704];
      10'd523 : out <= in [16767:16736];
      10'd524 : out <= in [16799:16768];
      10'd525 : out <= in [16831:16800];
      10'd526 : out <= in [16863:16832];
      10'd527 : out <= in [16895:16864];
      10'd528 : out <= in [16927:16896];
      10'd529 : out <= in [16959:16928];
      10'd530 : out <= in [16991:16960];
      10'd531 : out <= in [17023:16992];
      10'd532 : out <= in [17055:17024];
      10'd533 : out <= in [17087:17056];
      10'd534 : out <= in [17119:17088];
      10'd535 : out <= in [17151:17120];
      10'd536 : out <= in [17183:17152];
      10'd537 : out <= in [17215:17184];
      10'd538 : out <= in [17247:17216];
      10'd539 : out <= in [17279:17248];
      10'd540 : out <= in [17311:17280];
      10'd541 : out <= in [17343:17312];
      10'd542 : out <= in [17375:17344];
      10'd543 : out <= in [17407:17376];
      10'd544 : out <= in [17439:17408];
      10'd545 : out <= in [17471:17440];
      10'd546 : out <= in [17503:17472];
      10'd547 : out <= in [17535:17504];
      10'd548 : out <= in [17567:17536];
      10'd549 : out <= in [17599:17568];
      10'd550 : out <= in [17631:17600];
      10'd551 : out <= in [17663:17632];
      10'd552 : out <= in [17695:17664];
      10'd553 : out <= in [17727:17696];
      10'd554 : out <= in [17759:17728];
      10'd555 : out <= in [17791:17760];
      10'd556 : out <= in [17823:17792];
      10'd557 : out <= in [17855:17824];
      10'd558 : out <= in [17887:17856];
      10'd559 : out <= in [17919:17888];
      10'd560 : out <= in [17951:17920];
      10'd561 : out <= in [17983:17952];
      10'd562 : out <= in [18015:17984];
      10'd563 : out <= in [18047:18016];
      10'd564 : out <= in [18079:18048];
      10'd565 : out <= in [18111:18080];
      10'd566 : out <= in [18143:18112];
      10'd567 : out <= in [18175:18144];
      10'd568 : out <= in [18207:18176];
      10'd569 : out <= in [18239:18208];
      10'd570 : out <= in [18271:18240];
      10'd571 : out <= in [18303:18272];
      10'd572 : out <= in [18335:18304];
      10'd573 : out <= in [18367:18336];
      10'd574 : out <= in [18399:18368];
      10'd575 : out <= in [18431:18400];
      10'd576 : out <= in [18463:18432];
      10'd577 : out <= in [18495:18464];
      10'd578 : out <= in [18527:18496];
      10'd579 : out <= in [18559:18528];
      10'd580 : out <= in [18591:18560];
      10'd581 : out <= in [18623:18592];
      10'd582 : out <= in [18655:18624];
      10'd583 : out <= in [18687:18656];
      10'd584 : out <= in [18719:18688];
      10'd585 : out <= in [18751:18720];
      10'd586 : out <= in [18783:18752];
      10'd587 : out <= in [18815:18784];
      10'd588 : out <= in [18847:18816];
      10'd589 : out <= in [18879:18848];
      10'd590 : out <= in [18911:18880];
      10'd591 : out <= in [18943:18912];
      10'd592 : out <= in [18975:18944];
      10'd593 : out <= in [19007:18976];
      10'd594 : out <= in [19039:19008];
      10'd595 : out <= in [19071:19040];
      10'd596 : out <= in [19103:19072];
      10'd597 : out <= in [19135:19104];
      10'd598 : out <= in [19167:19136];
      10'd599 : out <= in [19199:19168];
      10'd600 : out <= in [19231:19200];
      10'd601 : out <= in [19263:19232];
      10'd602 : out <= in [19295:19264];
      10'd603 : out <= in [19327:19296];
      10'd604 : out <= in [19359:19328];
      10'd605 : out <= in [19391:19360];
      10'd606 : out <= in [19423:19392];
      10'd607 : out <= in [19455:19424];
      10'd608 : out <= in [19487:19456];
      10'd609 : out <= in [19519:19488];
      10'd610 : out <= in [19551:19520];
      10'd611 : out <= in [19583:19552];
      10'd612 : out <= in [19615:19584];
      10'd613 : out <= in [19647:19616];
      10'd614 : out <= in [19679:19648];
      10'd615 : out <= in [19711:19680];
      10'd616 : out <= in [19743:19712];
      10'd617 : out <= in [19775:19744];
      10'd618 : out <= in [19807:19776];
      10'd619 : out <= in [19839:19808];
      10'd620 : out <= in [19871:19840];
      10'd621 : out <= in [19903:19872];
      10'd622 : out <= in [19935:19904];
      10'd623 : out <= in [19967:19936];
      10'd624 : out <= in [19999:19968];
      10'd625 : out <= in [20031:20000];
      10'd626 : out <= in [20063:20032];
      10'd627 : out <= in [20095:20064];
      10'd628 : out <= in [20127:20096];
      10'd629 : out <= in [20159:20128];
      10'd630 : out <= in [20191:20160];
      10'd631 : out <= in [20223:20192];
      10'd632 : out <= in [20255:20224];
      10'd633 : out <= in [20287:20256];
      10'd634 : out <= in [20319:20288];
      10'd635 : out <= in [20351:20320];
      10'd636 : out <= in [20383:20352];
      10'd637 : out <= in [20415:20384];
      10'd638 : out <= in [20447:20416];
      10'd639 : out <= in [20479:20448];
      10'd640 : out <= in [20511:20480];
      10'd641 : out <= in [20543:20512];
      10'd642 : out <= in [20575:20544];
      10'd643 : out <= in [20607:20576];
      10'd644 : out <= in [20639:20608];
      10'd645 : out <= in [20671:20640];
      10'd646 : out <= in [20703:20672];
      10'd647 : out <= in [20735:20704];
      10'd648 : out <= in [20767:20736];
      10'd649 : out <= in [20799:20768];
      10'd650 : out <= in [20831:20800];
      10'd651 : out <= in [20863:20832];
      10'd652 : out <= in [20895:20864];
      10'd653 : out <= in [20927:20896];
      10'd654 : out <= in [20959:20928];
      10'd655 : out <= in [20991:20960];
      10'd656 : out <= in [21023:20992];
      10'd657 : out <= in [21055:21024];
      10'd658 : out <= in [21087:21056];
      10'd659 : out <= in [21119:21088];
      10'd660 : out <= in [21151:21120];
      10'd661 : out <= in [21183:21152];
      10'd662 : out <= in [21215:21184];
      10'd663 : out <= in [21247:21216];
      10'd664 : out <= in [21279:21248];
      10'd665 : out <= in [21311:21280];
      10'd666 : out <= in [21343:21312];
      10'd667 : out <= in [21375:21344];
      10'd668 : out <= in [21407:21376];
      10'd669 : out <= in [21439:21408];
      10'd670 : out <= in [21471:21440];
      10'd671 : out <= in [21503:21472];
      10'd672 : out <= in [21535:21504];
      10'd673 : out <= in [21567:21536];
      10'd674 : out <= in [21599:21568];
      10'd675 : out <= in [21631:21600];
      10'd676 : out <= in [21663:21632];
      10'd677 : out <= in [21695:21664];
      10'd678 : out <= in [21727:21696];
      10'd679 : out <= in [21759:21728];
      10'd680 : out <= in [21791:21760];
      10'd681 : out <= in [21823:21792];
      10'd682 : out <= in [21855:21824];
      10'd683 : out <= in [21887:21856];
      10'd684 : out <= in [21919:21888];
      10'd685 : out <= in [21951:21920];
      10'd686 : out <= in [21983:21952];
      10'd687 : out <= in [22015:21984];
      10'd688 : out <= in [22047:22016];
      10'd689 : out <= in [22079:22048];
      10'd690 : out <= in [22111:22080];
      10'd691 : out <= in [22143:22112];
      10'd692 : out <= in [22175:22144];
      10'd693 : out <= in [22207:22176];
      10'd694 : out <= in [22239:22208];
      10'd695 : out <= in [22271:22240];
      10'd696 : out <= in [22303:22272];
      10'd697 : out <= in [22335:22304];
      10'd698 : out <= in [22367:22336];
      10'd699 : out <= in [22399:22368];
      10'd700 : out <= in [22431:22400];
      10'd701 : out <= in [22463:22432];
      10'd702 : out <= in [22495:22464];
      10'd703 : out <= in [22527:22496];
      10'd704 : out <= in [22559:22528];
      10'd705 : out <= in [22591:22560];
      10'd706 : out <= in [22623:22592];
      10'd707 : out <= in [22655:22624];
      10'd708 : out <= in [22687:22656];
      10'd709 : out <= in [22719:22688];
      10'd710 : out <= in [22751:22720];
      10'd711 : out <= in [22783:22752];
      10'd712 : out <= in [22815:22784];
      10'd713 : out <= in [22847:22816];
      10'd714 : out <= in [22879:22848];
      10'd715 : out <= in [22911:22880];
      10'd716 : out <= in [22943:22912];
      10'd717 : out <= in [22975:22944];
      10'd718 : out <= in [23007:22976];
      10'd719 : out <= in [23039:23008];
      10'd720 : out <= in [23071:23040];
      10'd721 : out <= in [23103:23072];
      10'd722 : out <= in [23135:23104];
      10'd723 : out <= in [23167:23136];
      10'd724 : out <= in [23199:23168];
      10'd725 : out <= in [23231:23200];
      10'd726 : out <= in [23263:23232];
      10'd727 : out <= in [23295:23264];
      10'd728 : out <= in [23327:23296];
      10'd729 : out <= in [23359:23328];
      10'd730 : out <= in [23391:23360];
      10'd731 : out <= in [23423:23392];
      10'd732 : out <= in [23455:23424];
      10'd733 : out <= in [23487:23456];
      10'd734 : out <= in [23519:23488];
      10'd735 : out <= in [23551:23520];
      10'd736 : out <= in [23583:23552];
      10'd737 : out <= in [23615:23584];
      10'd738 : out <= in [23647:23616];
      10'd739 : out <= in [23679:23648];
      10'd740 : out <= in [23711:23680];
      10'd741 : out <= in [23743:23712];
      10'd742 : out <= in [23775:23744];
      10'd743 : out <= in [23807:23776];
      10'd744 : out <= in [23839:23808];
      10'd745 : out <= in [23871:23840];
      10'd746 : out <= in [23903:23872];
      10'd747 : out <= in [23935:23904];
      10'd748 : out <= in [23967:23936];
      10'd749 : out <= in [23999:23968];
      10'd750 : out <= in [24031:24000];
      10'd751 : out <= in [24063:24032];
      10'd752 : out <= in [24095:24064];
      10'd753 : out <= in [24127:24096];
      10'd754 : out <= in [24159:24128];
      10'd755 : out <= in [24191:24160];
      10'd756 : out <= in [24223:24192];
      10'd757 : out <= in [24255:24224];
      10'd758 : out <= in [24287:24256];
      10'd759 : out <= in [24319:24288];
      10'd760 : out <= in [24351:24320];
      10'd761 : out <= in [24383:24352];
      10'd762 : out <= in [24415:24384];
      10'd763 : out <= in [24447:24416];
      10'd764 : out <= in [24479:24448];
      10'd765 : out <= in [24511:24480];
      10'd766 : out <= in [24543:24512];
      10'd767 : out <= in [24575:24544];
      10'd768 : out <= in [24607:24576];
      10'd769 : out <= in [24639:24608];
      10'd770 : out <= in [24671:24640];
      10'd771 : out <= in [24703:24672];
      10'd772 : out <= in [24735:24704];
      10'd773 : out <= in [24767:24736];
      10'd774 : out <= in [24799:24768];
      10'd775 : out <= in [24831:24800];
      10'd776 : out <= in [24863:24832];
      10'd777 : out <= in [24895:24864];
      10'd778 : out <= in [24927:24896];
      10'd779 : out <= in [24959:24928];
      10'd780 : out <= in [24991:24960];
      10'd781 : out <= in [25023:24992];
      10'd782 : out <= in [25055:25024];
      10'd783 : out <= in [25087:25056];
      10'd784 : out <= in [25119:25088];
      10'd785 : out <= in [25151:25120];
      10'd786 : out <= in [25183:25152];
      10'd787 : out <= in [25215:25184];
      10'd788 : out <= in [25247:25216];
      10'd789 : out <= in [25279:25248];
      10'd790 : out <= in [25311:25280];
      10'd791 : out <= in [25343:25312];
      10'd792 : out <= in [25375:25344];
      10'd793 : out <= in [25407:25376];
      10'd794 : out <= in [25439:25408];
      10'd795 : out <= in [25471:25440];
      10'd796 : out <= in [25503:25472];
      10'd797 : out <= in [25535:25504];
      10'd798 : out <= in [25567:25536];
      10'd799 : out <= in [25599:25568];
      10'd800 : out <= in [25631:25600];
      10'd801 : out <= in [25663:25632];
      10'd802 : out <= in [25695:25664];
      10'd803 : out <= in [25727:25696];
      10'd804 : out <= in [25759:25728];
      10'd805 : out <= in [25791:25760];
      10'd806 : out <= in [25823:25792];
      10'd807 : out <= in [25855:25824];
      10'd808 : out <= in [25887:25856];
      10'd809 : out <= in [25919:25888];
      10'd810 : out <= in [25951:25920];
      10'd811 : out <= in [25983:25952];
      10'd812 : out <= in [26015:25984];
      10'd813 : out <= in [26047:26016];
      10'd814 : out <= in [26079:26048];
      10'd815 : out <= in [26111:26080];
      10'd816 : out <= in [26143:26112];
      10'd817 : out <= in [26175:26144];
      10'd818 : out <= in [26207:26176];
      10'd819 : out <= in [26239:26208];
      10'd820 : out <= in [26271:26240];
      10'd821 : out <= in [26303:26272];
      10'd822 : out <= in [26335:26304];
      10'd823 : out <= in [26367:26336];
      10'd824 : out <= in [26399:26368];
      10'd825 : out <= in [26431:26400];
      10'd826 : out <= in [26463:26432];
      10'd827 : out <= in [26495:26464];
      10'd828 : out <= in [26527:26496];
      10'd829 : out <= in [26559:26528];
      10'd830 : out <= in [26591:26560];
      10'd831 : out <= in [26623:26592];
      10'd832 : out <= in [26655:26624];
      10'd833 : out <= in [26687:26656];
      10'd834 : out <= in [26719:26688];
      10'd835 : out <= in [26751:26720];
      10'd836 : out <= in [26783:26752];
      10'd837 : out <= in [26815:26784];
      10'd838 : out <= in [26847:26816];
      10'd839 : out <= in [26879:26848];
      10'd840 : out <= in [26911:26880];
      10'd841 : out <= in [26943:26912];
      10'd842 : out <= in [26975:26944];
      10'd843 : out <= in [27007:26976];
      10'd844 : out <= in [27039:27008];
      10'd845 : out <= in [27071:27040];
      10'd846 : out <= in [27103:27072];
      10'd847 : out <= in [27135:27104];
      10'd848 : out <= in [27167:27136];
      10'd849 : out <= in [27199:27168];
      10'd850 : out <= in [27231:27200];
      10'd851 : out <= in [27263:27232];
      10'd852 : out <= in [27295:27264];
      10'd853 : out <= in [27327:27296];
      10'd854 : out <= in [27359:27328];
      10'd855 : out <= in [27391:27360];
      10'd856 : out <= in [27423:27392];
      10'd857 : out <= in [27455:27424];
      10'd858 : out <= in [27487:27456];
      10'd859 : out <= in [27519:27488];
      10'd860 : out <= in [27551:27520];
      10'd861 : out <= in [27583:27552];
      10'd862 : out <= in [27615:27584];
      10'd863 : out <= in [27647:27616];
      10'd864 : out <= in [27679:27648];
      10'd865 : out <= in [27711:27680];
      10'd866 : out <= in [27743:27712];
      10'd867 : out <= in [27775:27744];
      10'd868 : out <= in [27807:27776];
      10'd869 : out <= in [27839:27808];
      10'd870 : out <= in [27871:27840];
      10'd871 : out <= in [27903:27872];
      10'd872 : out <= in [27935:27904];
      10'd873 : out <= in [27967:27936];
      10'd874 : out <= in [27999:27968];
      10'd875 : out <= in [28031:28000];
      10'd876 : out <= in [28063:28032];
      10'd877 : out <= in [28095:28064];
      10'd878 : out <= in [28127:28096];
      10'd879 : out <= in [28159:28128];
      10'd880 : out <= in [28191:28160];
      10'd881 : out <= in [28223:28192];
      10'd882 : out <= in [28255:28224];
      10'd883 : out <= in [28287:28256];
      10'd884 : out <= in [28319:28288];
      10'd885 : out <= in [28351:28320];
      10'd886 : out <= in [28383:28352];
      10'd887 : out <= in [28415:28384];
      10'd888 : out <= in [28447:28416];
      10'd889 : out <= in [28479:28448];
      10'd890 : out <= in [28511:28480];
      10'd891 : out <= in [28543:28512];
      10'd892 : out <= in [28575:28544];
      10'd893 : out <= in [28607:28576];
      10'd894 : out <= in [28639:28608];
      10'd895 : out <= in [28671:28640];
      10'd896 : out <= in [28703:28672];
      10'd897 : out <= in [28735:28704];
      10'd898 : out <= in [28767:28736];
      10'd899 : out <= in [28799:28768];
      10'd900 : out <= in [28831:28800];
      10'd901 : out <= in [28863:28832];
      10'd902 : out <= in [28895:28864];
      10'd903 : out <= in [28927:28896];
      10'd904 : out <= in [28959:28928];
      10'd905 : out <= in [28991:28960];
      10'd906 : out <= in [29023:28992];
      10'd907 : out <= in [29055:29024];
      10'd908 : out <= in [29087:29056];
      10'd909 : out <= in [29119:29088];
      10'd910 : out <= in [29151:29120];
      10'd911 : out <= in [29183:29152];
      10'd912 : out <= in [29215:29184];
      10'd913 : out <= in [29247:29216];
      10'd914 : out <= in [29279:29248];
      10'd915 : out <= in [29311:29280];
      10'd916 : out <= in [29343:29312];
      10'd917 : out <= in [29375:29344];
      10'd918 : out <= in [29407:29376];
      10'd919 : out <= in [29439:29408];
      10'd920 : out <= in [29471:29440];
      10'd921 : out <= in [29503:29472];
      10'd922 : out <= in [29535:29504];
      10'd923 : out <= in [29567:29536];
      10'd924 : out <= in [29599:29568];
      10'd925 : out <= in [29631:29600];
      10'd926 : out <= in [29663:29632];
      10'd927 : out <= in [29695:29664];
      10'd928 : out <= in [29727:29696];
      10'd929 : out <= in [29759:29728];
      10'd930 : out <= in [29791:29760];
      10'd931 : out <= in [29823:29792];
      10'd932 : out <= in [29855:29824];
      10'd933 : out <= in [29887:29856];
      10'd934 : out <= in [29919:29888];
      10'd935 : out <= in [29951:29920];
      10'd936 : out <= in [29983:29952];
      10'd937 : out <= in [30015:29984];
      10'd938 : out <= in [30047:30016];
      10'd939 : out <= in [30079:30048];
      10'd940 : out <= in [30111:30080];
      10'd941 : out <= in [30143:30112];
      10'd942 : out <= in [30175:30144];
      10'd943 : out <= in [30207:30176];
      10'd944 : out <= in [30239:30208];
      10'd945 : out <= in [30271:30240];
      10'd946 : out <= in [30303:30272];
      10'd947 : out <= in [30335:30304];
      10'd948 : out <= in [30367:30336];
      10'd949 : out <= in [30399:30368];
      10'd950 : out <= in [30431:30400];
      10'd951 : out <= in [30463:30432];
      10'd952 : out <= in [30495:30464];
      10'd953 : out <= in [30527:30496];
      10'd954 : out <= in [30559:30528];
      10'd955 : out <= in [30591:30560];
      10'd956 : out <= in [30623:30592];
      10'd957 : out <= in [30655:30624];
      10'd958 : out <= in [30687:30656];
      10'd959 : out <= in [30719:30688];
      10'd960 : out <= in [30751:30720];
      10'd961 : out <= in [30783:30752];
      10'd962 : out <= in [30815:30784];
      10'd963 : out <= in [30847:30816];
      10'd964 : out <= in [30879:30848];
      10'd965 : out <= in [30911:30880];
      10'd966 : out <= in [30943:30912];
      10'd967 : out <= in [30975:30944];
      10'd968 : out <= in [31007:30976];
      10'd969 : out <= in [31039:31008];
      10'd970 : out <= in [31071:31040];
      10'd971 : out <= in [31103:31072];
      10'd972 : out <= in [31135:31104];
      10'd973 : out <= in [31167:31136];
      10'd974 : out <= in [31199:31168];
      10'd975 : out <= in [31231:31200];
      10'd976 : out <= in [31263:31232];
      10'd977 : out <= in [31295:31264];
      10'd978 : out <= in [31327:31296];
      10'd979 : out <= in [31359:31328];
      10'd980 : out <= in [31391:31360];
      10'd981 : out <= in [31423:31392];
      10'd982 : out <= in [31455:31424];
      10'd983 : out <= in [31487:31456];
      10'd984 : out <= in [31519:31488];
      10'd985 : out <= in [31551:31520];
      10'd986 : out <= in [31583:31552];
      10'd987 : out <= in [31615:31584];
      10'd988 : out <= in [31647:31616];
      10'd989 : out <= in [31679:31648];
      10'd990 : out <= in [31711:31680];
      10'd991 : out <= in [31743:31712];
      10'd992 : out <= in [31775:31744];
      10'd993 : out <= in [31807:31776];
      10'd994 : out <= in [31839:31808];
      10'd995 : out <= in [31871:31840];
      10'd996 : out <= in [31903:31872];
      10'd997 : out <= in [31935:31904];
      10'd998 : out <= in [31967:31936];
      10'd999 : out <= in [31999:31968];
      10'd1000 : out <= in [32031:32000];
      10'd1001 : out <= in [32063:32032];
      10'd1002 : out <= in [32095:32064];
      10'd1003 : out <= in [32127:32096];
      10'd1004 : out <= in [32159:32128];
      10'd1005 : out <= in [32191:32160];
      10'd1006 : out <= in [32223:32192];
      10'd1007 : out <= in [32255:32224];
      10'd1008 : out <= in [32287:32256];
      10'd1009 : out <= in [32319:32288];
      10'd1010 : out <= in [32351:32320];
      10'd1011 : out <= in [32383:32352];
      10'd1012 : out <= in [32415:32384];
      10'd1013 : out <= in [32447:32416];
      10'd1014 : out <= in [32479:32448];
      10'd1015 : out <= in [32511:32480];
      10'd1016 : out <= in [32543:32512];
      10'd1017 : out <= in [32575:32544];
      10'd1018 : out <= in [32607:32576];
      10'd1019 : out <= in [32639:32608];
      10'd1020 : out <= in [32671:32640];
      10'd1021 : out <= in [32703:32672];
      10'd1022 : out <= in [32735:32704];
      10'd1023 : out <= in [32767:32736];
      default: out <= 32'hxxxxxxxx;
    endcase
  end
endmodule

