module ready_bits_demux(
    in,
    addr,
    out,
    en
);

parameter TOTAL_INFO_LENGTH = `ISSUE_GPR_RD_BITS_LENGTH;

input [TOTAL_INFO_LENGTH-1:0] in;
input [`WF_ID_LENGTH-1:0] addr;
output [TOTAL_INFO_LENGTH*`WF_PER_CU-1:0] out;
reg [TOTAL_INFO_LENGTH*`WF_PER_CU-1:0] out;
input en;

always @(addr or in or en) begin
    out <= {(TOTAL_INFO_LENGTH*`WF_PER_CU-1){1'b0}};
    case(addr)
// %%start_veriperl
// my $i;
// for($i=0; $i<40; $i=$i+1)
// {
//   print "        6'd$i : out[TOTAL_INFO_LENGTH*$i+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*$i] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;\n";
// }
// %%stop_veriperl
        6'd0 : out[TOTAL_INFO_LENGTH*0+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*0] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd1 : out[TOTAL_INFO_LENGTH*1+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*1] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd2 : out[TOTAL_INFO_LENGTH*2+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*2] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd3 : out[TOTAL_INFO_LENGTH*3+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*3] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd4 : out[TOTAL_INFO_LENGTH*4+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*4] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd5 : out[TOTAL_INFO_LENGTH*5+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*5] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd6 : out[TOTAL_INFO_LENGTH*6+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*6] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd7 : out[TOTAL_INFO_LENGTH*7+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*7] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd8 : out[TOTAL_INFO_LENGTH*8+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*8] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd9 : out[TOTAL_INFO_LENGTH*9+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*9] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd10 : out[TOTAL_INFO_LENGTH*10+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*10] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd11 : out[TOTAL_INFO_LENGTH*11+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*11] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd12 : out[TOTAL_INFO_LENGTH*12+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*12] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd13 : out[TOTAL_INFO_LENGTH*13+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*13] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd14 : out[TOTAL_INFO_LENGTH*14+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*14] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd15 : out[TOTAL_INFO_LENGTH*15+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*15] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd16 : out[TOTAL_INFO_LENGTH*16+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*16] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd17 : out[TOTAL_INFO_LENGTH*17+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*17] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd18 : out[TOTAL_INFO_LENGTH*18+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*18] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd19 : out[TOTAL_INFO_LENGTH*19+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*19] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd20 : out[TOTAL_INFO_LENGTH*20+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*20] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd21 : out[TOTAL_INFO_LENGTH*21+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*21] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd22 : out[TOTAL_INFO_LENGTH*22+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*22] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd23 : out[TOTAL_INFO_LENGTH*23+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*23] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd24 : out[TOTAL_INFO_LENGTH*24+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*24] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd25 : out[TOTAL_INFO_LENGTH*25+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*25] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd26 : out[TOTAL_INFO_LENGTH*26+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*26] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd27 : out[TOTAL_INFO_LENGTH*27+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*27] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd28 : out[TOTAL_INFO_LENGTH*28+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*28] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd29 : out[TOTAL_INFO_LENGTH*29+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*29] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd30 : out[TOTAL_INFO_LENGTH*30+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*30] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd31 : out[TOTAL_INFO_LENGTH*31+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*31] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd32 : out[TOTAL_INFO_LENGTH*32+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*32] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd33 : out[TOTAL_INFO_LENGTH*33+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*33] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd34 : out[TOTAL_INFO_LENGTH*34+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*34] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd35 : out[TOTAL_INFO_LENGTH*35+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*35] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd36 : out[TOTAL_INFO_LENGTH*36+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*36] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd37 : out[TOTAL_INFO_LENGTH*37+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*37] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd38 : out[TOTAL_INFO_LENGTH*38+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*38] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
        6'd39 : out[TOTAL_INFO_LENGTH*39+(TOTAL_INFO_LENGTH-1):TOTAL_INFO_LENGTH*39] <= (en)? in: {TOTAL_INFO_LENGTH{1'b0}} ;
    endcase
end

endmodule
