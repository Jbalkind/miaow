module decoder_9_to_512 (out,in);
  output [511:0] out;
  input [8:0] in;
// %%start_veriperl
// my $i;
// for($i=0; $i<512; $i=$i+1)
// {
//   print "  assign out[$i] = (in == 9'd$i) ? 1'b1 : 1'b0;\n";
// }
// %%stop_veriperl
  assign out[0] = (in == 9'd0) ? 1'b1 : 1'b0;
  assign out[1] = (in == 9'd1) ? 1'b1 : 1'b0;
  assign out[2] = (in == 9'd2) ? 1'b1 : 1'b0;
  assign out[3] = (in == 9'd3) ? 1'b1 : 1'b0;
  assign out[4] = (in == 9'd4) ? 1'b1 : 1'b0;
  assign out[5] = (in == 9'd5) ? 1'b1 : 1'b0;
  assign out[6] = (in == 9'd6) ? 1'b1 : 1'b0;
  assign out[7] = (in == 9'd7) ? 1'b1 : 1'b0;
  assign out[8] = (in == 9'd8) ? 1'b1 : 1'b0;
  assign out[9] = (in == 9'd9) ? 1'b1 : 1'b0;
  assign out[10] = (in == 9'd10) ? 1'b1 : 1'b0;
  assign out[11] = (in == 9'd11) ? 1'b1 : 1'b0;
  assign out[12] = (in == 9'd12) ? 1'b1 : 1'b0;
  assign out[13] = (in == 9'd13) ? 1'b1 : 1'b0;
  assign out[14] = (in == 9'd14) ? 1'b1 : 1'b0;
  assign out[15] = (in == 9'd15) ? 1'b1 : 1'b0;
  assign out[16] = (in == 9'd16) ? 1'b1 : 1'b0;
  assign out[17] = (in == 9'd17) ? 1'b1 : 1'b0;
  assign out[18] = (in == 9'd18) ? 1'b1 : 1'b0;
  assign out[19] = (in == 9'd19) ? 1'b1 : 1'b0;
  assign out[20] = (in == 9'd20) ? 1'b1 : 1'b0;
  assign out[21] = (in == 9'd21) ? 1'b1 : 1'b0;
  assign out[22] = (in == 9'd22) ? 1'b1 : 1'b0;
  assign out[23] = (in == 9'd23) ? 1'b1 : 1'b0;
  assign out[24] = (in == 9'd24) ? 1'b1 : 1'b0;
  assign out[25] = (in == 9'd25) ? 1'b1 : 1'b0;
  assign out[26] = (in == 9'd26) ? 1'b1 : 1'b0;
  assign out[27] = (in == 9'd27) ? 1'b1 : 1'b0;
  assign out[28] = (in == 9'd28) ? 1'b1 : 1'b0;
  assign out[29] = (in == 9'd29) ? 1'b1 : 1'b0;
  assign out[30] = (in == 9'd30) ? 1'b1 : 1'b0;
  assign out[31] = (in == 9'd31) ? 1'b1 : 1'b0;
  assign out[32] = (in == 9'd32) ? 1'b1 : 1'b0;
  assign out[33] = (in == 9'd33) ? 1'b1 : 1'b0;
  assign out[34] = (in == 9'd34) ? 1'b1 : 1'b0;
  assign out[35] = (in == 9'd35) ? 1'b1 : 1'b0;
  assign out[36] = (in == 9'd36) ? 1'b1 : 1'b0;
  assign out[37] = (in == 9'd37) ? 1'b1 : 1'b0;
  assign out[38] = (in == 9'd38) ? 1'b1 : 1'b0;
  assign out[39] = (in == 9'd39) ? 1'b1 : 1'b0;
  assign out[40] = (in == 9'd40) ? 1'b1 : 1'b0;
  assign out[41] = (in == 9'd41) ? 1'b1 : 1'b0;
  assign out[42] = (in == 9'd42) ? 1'b1 : 1'b0;
  assign out[43] = (in == 9'd43) ? 1'b1 : 1'b0;
  assign out[44] = (in == 9'd44) ? 1'b1 : 1'b0;
  assign out[45] = (in == 9'd45) ? 1'b1 : 1'b0;
  assign out[46] = (in == 9'd46) ? 1'b1 : 1'b0;
  assign out[47] = (in == 9'd47) ? 1'b1 : 1'b0;
  assign out[48] = (in == 9'd48) ? 1'b1 : 1'b0;
  assign out[49] = (in == 9'd49) ? 1'b1 : 1'b0;
  assign out[50] = (in == 9'd50) ? 1'b1 : 1'b0;
  assign out[51] = (in == 9'd51) ? 1'b1 : 1'b0;
  assign out[52] = (in == 9'd52) ? 1'b1 : 1'b0;
  assign out[53] = (in == 9'd53) ? 1'b1 : 1'b0;
  assign out[54] = (in == 9'd54) ? 1'b1 : 1'b0;
  assign out[55] = (in == 9'd55) ? 1'b1 : 1'b0;
  assign out[56] = (in == 9'd56) ? 1'b1 : 1'b0;
  assign out[57] = (in == 9'd57) ? 1'b1 : 1'b0;
  assign out[58] = (in == 9'd58) ? 1'b1 : 1'b0;
  assign out[59] = (in == 9'd59) ? 1'b1 : 1'b0;
  assign out[60] = (in == 9'd60) ? 1'b1 : 1'b0;
  assign out[61] = (in == 9'd61) ? 1'b1 : 1'b0;
  assign out[62] = (in == 9'd62) ? 1'b1 : 1'b0;
  assign out[63] = (in == 9'd63) ? 1'b1 : 1'b0;
  assign out[64] = (in == 9'd64) ? 1'b1 : 1'b0;
  assign out[65] = (in == 9'd65) ? 1'b1 : 1'b0;
  assign out[66] = (in == 9'd66) ? 1'b1 : 1'b0;
  assign out[67] = (in == 9'd67) ? 1'b1 : 1'b0;
  assign out[68] = (in == 9'd68) ? 1'b1 : 1'b0;
  assign out[69] = (in == 9'd69) ? 1'b1 : 1'b0;
  assign out[70] = (in == 9'd70) ? 1'b1 : 1'b0;
  assign out[71] = (in == 9'd71) ? 1'b1 : 1'b0;
  assign out[72] = (in == 9'd72) ? 1'b1 : 1'b0;
  assign out[73] = (in == 9'd73) ? 1'b1 : 1'b0;
  assign out[74] = (in == 9'd74) ? 1'b1 : 1'b0;
  assign out[75] = (in == 9'd75) ? 1'b1 : 1'b0;
  assign out[76] = (in == 9'd76) ? 1'b1 : 1'b0;
  assign out[77] = (in == 9'd77) ? 1'b1 : 1'b0;
  assign out[78] = (in == 9'd78) ? 1'b1 : 1'b0;
  assign out[79] = (in == 9'd79) ? 1'b1 : 1'b0;
  assign out[80] = (in == 9'd80) ? 1'b1 : 1'b0;
  assign out[81] = (in == 9'd81) ? 1'b1 : 1'b0;
  assign out[82] = (in == 9'd82) ? 1'b1 : 1'b0;
  assign out[83] = (in == 9'd83) ? 1'b1 : 1'b0;
  assign out[84] = (in == 9'd84) ? 1'b1 : 1'b0;
  assign out[85] = (in == 9'd85) ? 1'b1 : 1'b0;
  assign out[86] = (in == 9'd86) ? 1'b1 : 1'b0;
  assign out[87] = (in == 9'd87) ? 1'b1 : 1'b0;
  assign out[88] = (in == 9'd88) ? 1'b1 : 1'b0;
  assign out[89] = (in == 9'd89) ? 1'b1 : 1'b0;
  assign out[90] = (in == 9'd90) ? 1'b1 : 1'b0;
  assign out[91] = (in == 9'd91) ? 1'b1 : 1'b0;
  assign out[92] = (in == 9'd92) ? 1'b1 : 1'b0;
  assign out[93] = (in == 9'd93) ? 1'b1 : 1'b0;
  assign out[94] = (in == 9'd94) ? 1'b1 : 1'b0;
  assign out[95] = (in == 9'd95) ? 1'b1 : 1'b0;
  assign out[96] = (in == 9'd96) ? 1'b1 : 1'b0;
  assign out[97] = (in == 9'd97) ? 1'b1 : 1'b0;
  assign out[98] = (in == 9'd98) ? 1'b1 : 1'b0;
  assign out[99] = (in == 9'd99) ? 1'b1 : 1'b0;
  assign out[100] = (in == 9'd100) ? 1'b1 : 1'b0;
  assign out[101] = (in == 9'd101) ? 1'b1 : 1'b0;
  assign out[102] = (in == 9'd102) ? 1'b1 : 1'b0;
  assign out[103] = (in == 9'd103) ? 1'b1 : 1'b0;
  assign out[104] = (in == 9'd104) ? 1'b1 : 1'b0;
  assign out[105] = (in == 9'd105) ? 1'b1 : 1'b0;
  assign out[106] = (in == 9'd106) ? 1'b1 : 1'b0;
  assign out[107] = (in == 9'd107) ? 1'b1 : 1'b0;
  assign out[108] = (in == 9'd108) ? 1'b1 : 1'b0;
  assign out[109] = (in == 9'd109) ? 1'b1 : 1'b0;
  assign out[110] = (in == 9'd110) ? 1'b1 : 1'b0;
  assign out[111] = (in == 9'd111) ? 1'b1 : 1'b0;
  assign out[112] = (in == 9'd112) ? 1'b1 : 1'b0;
  assign out[113] = (in == 9'd113) ? 1'b1 : 1'b0;
  assign out[114] = (in == 9'd114) ? 1'b1 : 1'b0;
  assign out[115] = (in == 9'd115) ? 1'b1 : 1'b0;
  assign out[116] = (in == 9'd116) ? 1'b1 : 1'b0;
  assign out[117] = (in == 9'd117) ? 1'b1 : 1'b0;
  assign out[118] = (in == 9'd118) ? 1'b1 : 1'b0;
  assign out[119] = (in == 9'd119) ? 1'b1 : 1'b0;
  assign out[120] = (in == 9'd120) ? 1'b1 : 1'b0;
  assign out[121] = (in == 9'd121) ? 1'b1 : 1'b0;
  assign out[122] = (in == 9'd122) ? 1'b1 : 1'b0;
  assign out[123] = (in == 9'd123) ? 1'b1 : 1'b0;
  assign out[124] = (in == 9'd124) ? 1'b1 : 1'b0;
  assign out[125] = (in == 9'd125) ? 1'b1 : 1'b0;
  assign out[126] = (in == 9'd126) ? 1'b1 : 1'b0;
  assign out[127] = (in == 9'd127) ? 1'b1 : 1'b0;
  assign out[128] = (in == 9'd128) ? 1'b1 : 1'b0;
  assign out[129] = (in == 9'd129) ? 1'b1 : 1'b0;
  assign out[130] = (in == 9'd130) ? 1'b1 : 1'b0;
  assign out[131] = (in == 9'd131) ? 1'b1 : 1'b0;
  assign out[132] = (in == 9'd132) ? 1'b1 : 1'b0;
  assign out[133] = (in == 9'd133) ? 1'b1 : 1'b0;
  assign out[134] = (in == 9'd134) ? 1'b1 : 1'b0;
  assign out[135] = (in == 9'd135) ? 1'b1 : 1'b0;
  assign out[136] = (in == 9'd136) ? 1'b1 : 1'b0;
  assign out[137] = (in == 9'd137) ? 1'b1 : 1'b0;
  assign out[138] = (in == 9'd138) ? 1'b1 : 1'b0;
  assign out[139] = (in == 9'd139) ? 1'b1 : 1'b0;
  assign out[140] = (in == 9'd140) ? 1'b1 : 1'b0;
  assign out[141] = (in == 9'd141) ? 1'b1 : 1'b0;
  assign out[142] = (in == 9'd142) ? 1'b1 : 1'b0;
  assign out[143] = (in == 9'd143) ? 1'b1 : 1'b0;
  assign out[144] = (in == 9'd144) ? 1'b1 : 1'b0;
  assign out[145] = (in == 9'd145) ? 1'b1 : 1'b0;
  assign out[146] = (in == 9'd146) ? 1'b1 : 1'b0;
  assign out[147] = (in == 9'd147) ? 1'b1 : 1'b0;
  assign out[148] = (in == 9'd148) ? 1'b1 : 1'b0;
  assign out[149] = (in == 9'd149) ? 1'b1 : 1'b0;
  assign out[150] = (in == 9'd150) ? 1'b1 : 1'b0;
  assign out[151] = (in == 9'd151) ? 1'b1 : 1'b0;
  assign out[152] = (in == 9'd152) ? 1'b1 : 1'b0;
  assign out[153] = (in == 9'd153) ? 1'b1 : 1'b0;
  assign out[154] = (in == 9'd154) ? 1'b1 : 1'b0;
  assign out[155] = (in == 9'd155) ? 1'b1 : 1'b0;
  assign out[156] = (in == 9'd156) ? 1'b1 : 1'b0;
  assign out[157] = (in == 9'd157) ? 1'b1 : 1'b0;
  assign out[158] = (in == 9'd158) ? 1'b1 : 1'b0;
  assign out[159] = (in == 9'd159) ? 1'b1 : 1'b0;
  assign out[160] = (in == 9'd160) ? 1'b1 : 1'b0;
  assign out[161] = (in == 9'd161) ? 1'b1 : 1'b0;
  assign out[162] = (in == 9'd162) ? 1'b1 : 1'b0;
  assign out[163] = (in == 9'd163) ? 1'b1 : 1'b0;
  assign out[164] = (in == 9'd164) ? 1'b1 : 1'b0;
  assign out[165] = (in == 9'd165) ? 1'b1 : 1'b0;
  assign out[166] = (in == 9'd166) ? 1'b1 : 1'b0;
  assign out[167] = (in == 9'd167) ? 1'b1 : 1'b0;
  assign out[168] = (in == 9'd168) ? 1'b1 : 1'b0;
  assign out[169] = (in == 9'd169) ? 1'b1 : 1'b0;
  assign out[170] = (in == 9'd170) ? 1'b1 : 1'b0;
  assign out[171] = (in == 9'd171) ? 1'b1 : 1'b0;
  assign out[172] = (in == 9'd172) ? 1'b1 : 1'b0;
  assign out[173] = (in == 9'd173) ? 1'b1 : 1'b0;
  assign out[174] = (in == 9'd174) ? 1'b1 : 1'b0;
  assign out[175] = (in == 9'd175) ? 1'b1 : 1'b0;
  assign out[176] = (in == 9'd176) ? 1'b1 : 1'b0;
  assign out[177] = (in == 9'd177) ? 1'b1 : 1'b0;
  assign out[178] = (in == 9'd178) ? 1'b1 : 1'b0;
  assign out[179] = (in == 9'd179) ? 1'b1 : 1'b0;
  assign out[180] = (in == 9'd180) ? 1'b1 : 1'b0;
  assign out[181] = (in == 9'd181) ? 1'b1 : 1'b0;
  assign out[182] = (in == 9'd182) ? 1'b1 : 1'b0;
  assign out[183] = (in == 9'd183) ? 1'b1 : 1'b0;
  assign out[184] = (in == 9'd184) ? 1'b1 : 1'b0;
  assign out[185] = (in == 9'd185) ? 1'b1 : 1'b0;
  assign out[186] = (in == 9'd186) ? 1'b1 : 1'b0;
  assign out[187] = (in == 9'd187) ? 1'b1 : 1'b0;
  assign out[188] = (in == 9'd188) ? 1'b1 : 1'b0;
  assign out[189] = (in == 9'd189) ? 1'b1 : 1'b0;
  assign out[190] = (in == 9'd190) ? 1'b1 : 1'b0;
  assign out[191] = (in == 9'd191) ? 1'b1 : 1'b0;
  assign out[192] = (in == 9'd192) ? 1'b1 : 1'b0;
  assign out[193] = (in == 9'd193) ? 1'b1 : 1'b0;
  assign out[194] = (in == 9'd194) ? 1'b1 : 1'b0;
  assign out[195] = (in == 9'd195) ? 1'b1 : 1'b0;
  assign out[196] = (in == 9'd196) ? 1'b1 : 1'b0;
  assign out[197] = (in == 9'd197) ? 1'b1 : 1'b0;
  assign out[198] = (in == 9'd198) ? 1'b1 : 1'b0;
  assign out[199] = (in == 9'd199) ? 1'b1 : 1'b0;
  assign out[200] = (in == 9'd200) ? 1'b1 : 1'b0;
  assign out[201] = (in == 9'd201) ? 1'b1 : 1'b0;
  assign out[202] = (in == 9'd202) ? 1'b1 : 1'b0;
  assign out[203] = (in == 9'd203) ? 1'b1 : 1'b0;
  assign out[204] = (in == 9'd204) ? 1'b1 : 1'b0;
  assign out[205] = (in == 9'd205) ? 1'b1 : 1'b0;
  assign out[206] = (in == 9'd206) ? 1'b1 : 1'b0;
  assign out[207] = (in == 9'd207) ? 1'b1 : 1'b0;
  assign out[208] = (in == 9'd208) ? 1'b1 : 1'b0;
  assign out[209] = (in == 9'd209) ? 1'b1 : 1'b0;
  assign out[210] = (in == 9'd210) ? 1'b1 : 1'b0;
  assign out[211] = (in == 9'd211) ? 1'b1 : 1'b0;
  assign out[212] = (in == 9'd212) ? 1'b1 : 1'b0;
  assign out[213] = (in == 9'd213) ? 1'b1 : 1'b0;
  assign out[214] = (in == 9'd214) ? 1'b1 : 1'b0;
  assign out[215] = (in == 9'd215) ? 1'b1 : 1'b0;
  assign out[216] = (in == 9'd216) ? 1'b1 : 1'b0;
  assign out[217] = (in == 9'd217) ? 1'b1 : 1'b0;
  assign out[218] = (in == 9'd218) ? 1'b1 : 1'b0;
  assign out[219] = (in == 9'd219) ? 1'b1 : 1'b0;
  assign out[220] = (in == 9'd220) ? 1'b1 : 1'b0;
  assign out[221] = (in == 9'd221) ? 1'b1 : 1'b0;
  assign out[222] = (in == 9'd222) ? 1'b1 : 1'b0;
  assign out[223] = (in == 9'd223) ? 1'b1 : 1'b0;
  assign out[224] = (in == 9'd224) ? 1'b1 : 1'b0;
  assign out[225] = (in == 9'd225) ? 1'b1 : 1'b0;
  assign out[226] = (in == 9'd226) ? 1'b1 : 1'b0;
  assign out[227] = (in == 9'd227) ? 1'b1 : 1'b0;
  assign out[228] = (in == 9'd228) ? 1'b1 : 1'b0;
  assign out[229] = (in == 9'd229) ? 1'b1 : 1'b0;
  assign out[230] = (in == 9'd230) ? 1'b1 : 1'b0;
  assign out[231] = (in == 9'd231) ? 1'b1 : 1'b0;
  assign out[232] = (in == 9'd232) ? 1'b1 : 1'b0;
  assign out[233] = (in == 9'd233) ? 1'b1 : 1'b0;
  assign out[234] = (in == 9'd234) ? 1'b1 : 1'b0;
  assign out[235] = (in == 9'd235) ? 1'b1 : 1'b0;
  assign out[236] = (in == 9'd236) ? 1'b1 : 1'b0;
  assign out[237] = (in == 9'd237) ? 1'b1 : 1'b0;
  assign out[238] = (in == 9'd238) ? 1'b1 : 1'b0;
  assign out[239] = (in == 9'd239) ? 1'b1 : 1'b0;
  assign out[240] = (in == 9'd240) ? 1'b1 : 1'b0;
  assign out[241] = (in == 9'd241) ? 1'b1 : 1'b0;
  assign out[242] = (in == 9'd242) ? 1'b1 : 1'b0;
  assign out[243] = (in == 9'd243) ? 1'b1 : 1'b0;
  assign out[244] = (in == 9'd244) ? 1'b1 : 1'b0;
  assign out[245] = (in == 9'd245) ? 1'b1 : 1'b0;
  assign out[246] = (in == 9'd246) ? 1'b1 : 1'b0;
  assign out[247] = (in == 9'd247) ? 1'b1 : 1'b0;
  assign out[248] = (in == 9'd248) ? 1'b1 : 1'b0;
  assign out[249] = (in == 9'd249) ? 1'b1 : 1'b0;
  assign out[250] = (in == 9'd250) ? 1'b1 : 1'b0;
  assign out[251] = (in == 9'd251) ? 1'b1 : 1'b0;
  assign out[252] = (in == 9'd252) ? 1'b1 : 1'b0;
  assign out[253] = (in == 9'd253) ? 1'b1 : 1'b0;
  assign out[254] = (in == 9'd254) ? 1'b1 : 1'b0;
  assign out[255] = (in == 9'd255) ? 1'b1 : 1'b0;
  assign out[256] = (in == 9'd256) ? 1'b1 : 1'b0;
  assign out[257] = (in == 9'd257) ? 1'b1 : 1'b0;
  assign out[258] = (in == 9'd258) ? 1'b1 : 1'b0;
  assign out[259] = (in == 9'd259) ? 1'b1 : 1'b0;
  assign out[260] = (in == 9'd260) ? 1'b1 : 1'b0;
  assign out[261] = (in == 9'd261) ? 1'b1 : 1'b0;
  assign out[262] = (in == 9'd262) ? 1'b1 : 1'b0;
  assign out[263] = (in == 9'd263) ? 1'b1 : 1'b0;
  assign out[264] = (in == 9'd264) ? 1'b1 : 1'b0;
  assign out[265] = (in == 9'd265) ? 1'b1 : 1'b0;
  assign out[266] = (in == 9'd266) ? 1'b1 : 1'b0;
  assign out[267] = (in == 9'd267) ? 1'b1 : 1'b0;
  assign out[268] = (in == 9'd268) ? 1'b1 : 1'b0;
  assign out[269] = (in == 9'd269) ? 1'b1 : 1'b0;
  assign out[270] = (in == 9'd270) ? 1'b1 : 1'b0;
  assign out[271] = (in == 9'd271) ? 1'b1 : 1'b0;
  assign out[272] = (in == 9'd272) ? 1'b1 : 1'b0;
  assign out[273] = (in == 9'd273) ? 1'b1 : 1'b0;
  assign out[274] = (in == 9'd274) ? 1'b1 : 1'b0;
  assign out[275] = (in == 9'd275) ? 1'b1 : 1'b0;
  assign out[276] = (in == 9'd276) ? 1'b1 : 1'b0;
  assign out[277] = (in == 9'd277) ? 1'b1 : 1'b0;
  assign out[278] = (in == 9'd278) ? 1'b1 : 1'b0;
  assign out[279] = (in == 9'd279) ? 1'b1 : 1'b0;
  assign out[280] = (in == 9'd280) ? 1'b1 : 1'b0;
  assign out[281] = (in == 9'd281) ? 1'b1 : 1'b0;
  assign out[282] = (in == 9'd282) ? 1'b1 : 1'b0;
  assign out[283] = (in == 9'd283) ? 1'b1 : 1'b0;
  assign out[284] = (in == 9'd284) ? 1'b1 : 1'b0;
  assign out[285] = (in == 9'd285) ? 1'b1 : 1'b0;
  assign out[286] = (in == 9'd286) ? 1'b1 : 1'b0;
  assign out[287] = (in == 9'd287) ? 1'b1 : 1'b0;
  assign out[288] = (in == 9'd288) ? 1'b1 : 1'b0;
  assign out[289] = (in == 9'd289) ? 1'b1 : 1'b0;
  assign out[290] = (in == 9'd290) ? 1'b1 : 1'b0;
  assign out[291] = (in == 9'd291) ? 1'b1 : 1'b0;
  assign out[292] = (in == 9'd292) ? 1'b1 : 1'b0;
  assign out[293] = (in == 9'd293) ? 1'b1 : 1'b0;
  assign out[294] = (in == 9'd294) ? 1'b1 : 1'b0;
  assign out[295] = (in == 9'd295) ? 1'b1 : 1'b0;
  assign out[296] = (in == 9'd296) ? 1'b1 : 1'b0;
  assign out[297] = (in == 9'd297) ? 1'b1 : 1'b0;
  assign out[298] = (in == 9'd298) ? 1'b1 : 1'b0;
  assign out[299] = (in == 9'd299) ? 1'b1 : 1'b0;
  assign out[300] = (in == 9'd300) ? 1'b1 : 1'b0;
  assign out[301] = (in == 9'd301) ? 1'b1 : 1'b0;
  assign out[302] = (in == 9'd302) ? 1'b1 : 1'b0;
  assign out[303] = (in == 9'd303) ? 1'b1 : 1'b0;
  assign out[304] = (in == 9'd304) ? 1'b1 : 1'b0;
  assign out[305] = (in == 9'd305) ? 1'b1 : 1'b0;
  assign out[306] = (in == 9'd306) ? 1'b1 : 1'b0;
  assign out[307] = (in == 9'd307) ? 1'b1 : 1'b0;
  assign out[308] = (in == 9'd308) ? 1'b1 : 1'b0;
  assign out[309] = (in == 9'd309) ? 1'b1 : 1'b0;
  assign out[310] = (in == 9'd310) ? 1'b1 : 1'b0;
  assign out[311] = (in == 9'd311) ? 1'b1 : 1'b0;
  assign out[312] = (in == 9'd312) ? 1'b1 : 1'b0;
  assign out[313] = (in == 9'd313) ? 1'b1 : 1'b0;
  assign out[314] = (in == 9'd314) ? 1'b1 : 1'b0;
  assign out[315] = (in == 9'd315) ? 1'b1 : 1'b0;
  assign out[316] = (in == 9'd316) ? 1'b1 : 1'b0;
  assign out[317] = (in == 9'd317) ? 1'b1 : 1'b0;
  assign out[318] = (in == 9'd318) ? 1'b1 : 1'b0;
  assign out[319] = (in == 9'd319) ? 1'b1 : 1'b0;
  assign out[320] = (in == 9'd320) ? 1'b1 : 1'b0;
  assign out[321] = (in == 9'd321) ? 1'b1 : 1'b0;
  assign out[322] = (in == 9'd322) ? 1'b1 : 1'b0;
  assign out[323] = (in == 9'd323) ? 1'b1 : 1'b0;
  assign out[324] = (in == 9'd324) ? 1'b1 : 1'b0;
  assign out[325] = (in == 9'd325) ? 1'b1 : 1'b0;
  assign out[326] = (in == 9'd326) ? 1'b1 : 1'b0;
  assign out[327] = (in == 9'd327) ? 1'b1 : 1'b0;
  assign out[328] = (in == 9'd328) ? 1'b1 : 1'b0;
  assign out[329] = (in == 9'd329) ? 1'b1 : 1'b0;
  assign out[330] = (in == 9'd330) ? 1'b1 : 1'b0;
  assign out[331] = (in == 9'd331) ? 1'b1 : 1'b0;
  assign out[332] = (in == 9'd332) ? 1'b1 : 1'b0;
  assign out[333] = (in == 9'd333) ? 1'b1 : 1'b0;
  assign out[334] = (in == 9'd334) ? 1'b1 : 1'b0;
  assign out[335] = (in == 9'd335) ? 1'b1 : 1'b0;
  assign out[336] = (in == 9'd336) ? 1'b1 : 1'b0;
  assign out[337] = (in == 9'd337) ? 1'b1 : 1'b0;
  assign out[338] = (in == 9'd338) ? 1'b1 : 1'b0;
  assign out[339] = (in == 9'd339) ? 1'b1 : 1'b0;
  assign out[340] = (in == 9'd340) ? 1'b1 : 1'b0;
  assign out[341] = (in == 9'd341) ? 1'b1 : 1'b0;
  assign out[342] = (in == 9'd342) ? 1'b1 : 1'b0;
  assign out[343] = (in == 9'd343) ? 1'b1 : 1'b0;
  assign out[344] = (in == 9'd344) ? 1'b1 : 1'b0;
  assign out[345] = (in == 9'd345) ? 1'b1 : 1'b0;
  assign out[346] = (in == 9'd346) ? 1'b1 : 1'b0;
  assign out[347] = (in == 9'd347) ? 1'b1 : 1'b0;
  assign out[348] = (in == 9'd348) ? 1'b1 : 1'b0;
  assign out[349] = (in == 9'd349) ? 1'b1 : 1'b0;
  assign out[350] = (in == 9'd350) ? 1'b1 : 1'b0;
  assign out[351] = (in == 9'd351) ? 1'b1 : 1'b0;
  assign out[352] = (in == 9'd352) ? 1'b1 : 1'b0;
  assign out[353] = (in == 9'd353) ? 1'b1 : 1'b0;
  assign out[354] = (in == 9'd354) ? 1'b1 : 1'b0;
  assign out[355] = (in == 9'd355) ? 1'b1 : 1'b0;
  assign out[356] = (in == 9'd356) ? 1'b1 : 1'b0;
  assign out[357] = (in == 9'd357) ? 1'b1 : 1'b0;
  assign out[358] = (in == 9'd358) ? 1'b1 : 1'b0;
  assign out[359] = (in == 9'd359) ? 1'b1 : 1'b0;
  assign out[360] = (in == 9'd360) ? 1'b1 : 1'b0;
  assign out[361] = (in == 9'd361) ? 1'b1 : 1'b0;
  assign out[362] = (in == 9'd362) ? 1'b1 : 1'b0;
  assign out[363] = (in == 9'd363) ? 1'b1 : 1'b0;
  assign out[364] = (in == 9'd364) ? 1'b1 : 1'b0;
  assign out[365] = (in == 9'd365) ? 1'b1 : 1'b0;
  assign out[366] = (in == 9'd366) ? 1'b1 : 1'b0;
  assign out[367] = (in == 9'd367) ? 1'b1 : 1'b0;
  assign out[368] = (in == 9'd368) ? 1'b1 : 1'b0;
  assign out[369] = (in == 9'd369) ? 1'b1 : 1'b0;
  assign out[370] = (in == 9'd370) ? 1'b1 : 1'b0;
  assign out[371] = (in == 9'd371) ? 1'b1 : 1'b0;
  assign out[372] = (in == 9'd372) ? 1'b1 : 1'b0;
  assign out[373] = (in == 9'd373) ? 1'b1 : 1'b0;
  assign out[374] = (in == 9'd374) ? 1'b1 : 1'b0;
  assign out[375] = (in == 9'd375) ? 1'b1 : 1'b0;
  assign out[376] = (in == 9'd376) ? 1'b1 : 1'b0;
  assign out[377] = (in == 9'd377) ? 1'b1 : 1'b0;
  assign out[378] = (in == 9'd378) ? 1'b1 : 1'b0;
  assign out[379] = (in == 9'd379) ? 1'b1 : 1'b0;
  assign out[380] = (in == 9'd380) ? 1'b1 : 1'b0;
  assign out[381] = (in == 9'd381) ? 1'b1 : 1'b0;
  assign out[382] = (in == 9'd382) ? 1'b1 : 1'b0;
  assign out[383] = (in == 9'd383) ? 1'b1 : 1'b0;
  assign out[384] = (in == 9'd384) ? 1'b1 : 1'b0;
  assign out[385] = (in == 9'd385) ? 1'b1 : 1'b0;
  assign out[386] = (in == 9'd386) ? 1'b1 : 1'b0;
  assign out[387] = (in == 9'd387) ? 1'b1 : 1'b0;
  assign out[388] = (in == 9'd388) ? 1'b1 : 1'b0;
  assign out[389] = (in == 9'd389) ? 1'b1 : 1'b0;
  assign out[390] = (in == 9'd390) ? 1'b1 : 1'b0;
  assign out[391] = (in == 9'd391) ? 1'b1 : 1'b0;
  assign out[392] = (in == 9'd392) ? 1'b1 : 1'b0;
  assign out[393] = (in == 9'd393) ? 1'b1 : 1'b0;
  assign out[394] = (in == 9'd394) ? 1'b1 : 1'b0;
  assign out[395] = (in == 9'd395) ? 1'b1 : 1'b0;
  assign out[396] = (in == 9'd396) ? 1'b1 : 1'b0;
  assign out[397] = (in == 9'd397) ? 1'b1 : 1'b0;
  assign out[398] = (in == 9'd398) ? 1'b1 : 1'b0;
  assign out[399] = (in == 9'd399) ? 1'b1 : 1'b0;
  assign out[400] = (in == 9'd400) ? 1'b1 : 1'b0;
  assign out[401] = (in == 9'd401) ? 1'b1 : 1'b0;
  assign out[402] = (in == 9'd402) ? 1'b1 : 1'b0;
  assign out[403] = (in == 9'd403) ? 1'b1 : 1'b0;
  assign out[404] = (in == 9'd404) ? 1'b1 : 1'b0;
  assign out[405] = (in == 9'd405) ? 1'b1 : 1'b0;
  assign out[406] = (in == 9'd406) ? 1'b1 : 1'b0;
  assign out[407] = (in == 9'd407) ? 1'b1 : 1'b0;
  assign out[408] = (in == 9'd408) ? 1'b1 : 1'b0;
  assign out[409] = (in == 9'd409) ? 1'b1 : 1'b0;
  assign out[410] = (in == 9'd410) ? 1'b1 : 1'b0;
  assign out[411] = (in == 9'd411) ? 1'b1 : 1'b0;
  assign out[412] = (in == 9'd412) ? 1'b1 : 1'b0;
  assign out[413] = (in == 9'd413) ? 1'b1 : 1'b0;
  assign out[414] = (in == 9'd414) ? 1'b1 : 1'b0;
  assign out[415] = (in == 9'd415) ? 1'b1 : 1'b0;
  assign out[416] = (in == 9'd416) ? 1'b1 : 1'b0;
  assign out[417] = (in == 9'd417) ? 1'b1 : 1'b0;
  assign out[418] = (in == 9'd418) ? 1'b1 : 1'b0;
  assign out[419] = (in == 9'd419) ? 1'b1 : 1'b0;
  assign out[420] = (in == 9'd420) ? 1'b1 : 1'b0;
  assign out[421] = (in == 9'd421) ? 1'b1 : 1'b0;
  assign out[422] = (in == 9'd422) ? 1'b1 : 1'b0;
  assign out[423] = (in == 9'd423) ? 1'b1 : 1'b0;
  assign out[424] = (in == 9'd424) ? 1'b1 : 1'b0;
  assign out[425] = (in == 9'd425) ? 1'b1 : 1'b0;
  assign out[426] = (in == 9'd426) ? 1'b1 : 1'b0;
  assign out[427] = (in == 9'd427) ? 1'b1 : 1'b0;
  assign out[428] = (in == 9'd428) ? 1'b1 : 1'b0;
  assign out[429] = (in == 9'd429) ? 1'b1 : 1'b0;
  assign out[430] = (in == 9'd430) ? 1'b1 : 1'b0;
  assign out[431] = (in == 9'd431) ? 1'b1 : 1'b0;
  assign out[432] = (in == 9'd432) ? 1'b1 : 1'b0;
  assign out[433] = (in == 9'd433) ? 1'b1 : 1'b0;
  assign out[434] = (in == 9'd434) ? 1'b1 : 1'b0;
  assign out[435] = (in == 9'd435) ? 1'b1 : 1'b0;
  assign out[436] = (in == 9'd436) ? 1'b1 : 1'b0;
  assign out[437] = (in == 9'd437) ? 1'b1 : 1'b0;
  assign out[438] = (in == 9'd438) ? 1'b1 : 1'b0;
  assign out[439] = (in == 9'd439) ? 1'b1 : 1'b0;
  assign out[440] = (in == 9'd440) ? 1'b1 : 1'b0;
  assign out[441] = (in == 9'd441) ? 1'b1 : 1'b0;
  assign out[442] = (in == 9'd442) ? 1'b1 : 1'b0;
  assign out[443] = (in == 9'd443) ? 1'b1 : 1'b0;
  assign out[444] = (in == 9'd444) ? 1'b1 : 1'b0;
  assign out[445] = (in == 9'd445) ? 1'b1 : 1'b0;
  assign out[446] = (in == 9'd446) ? 1'b1 : 1'b0;
  assign out[447] = (in == 9'd447) ? 1'b1 : 1'b0;
  assign out[448] = (in == 9'd448) ? 1'b1 : 1'b0;
  assign out[449] = (in == 9'd449) ? 1'b1 : 1'b0;
  assign out[450] = (in == 9'd450) ? 1'b1 : 1'b0;
  assign out[451] = (in == 9'd451) ? 1'b1 : 1'b0;
  assign out[452] = (in == 9'd452) ? 1'b1 : 1'b0;
  assign out[453] = (in == 9'd453) ? 1'b1 : 1'b0;
  assign out[454] = (in == 9'd454) ? 1'b1 : 1'b0;
  assign out[455] = (in == 9'd455) ? 1'b1 : 1'b0;
  assign out[456] = (in == 9'd456) ? 1'b1 : 1'b0;
  assign out[457] = (in == 9'd457) ? 1'b1 : 1'b0;
  assign out[458] = (in == 9'd458) ? 1'b1 : 1'b0;
  assign out[459] = (in == 9'd459) ? 1'b1 : 1'b0;
  assign out[460] = (in == 9'd460) ? 1'b1 : 1'b0;
  assign out[461] = (in == 9'd461) ? 1'b1 : 1'b0;
  assign out[462] = (in == 9'd462) ? 1'b1 : 1'b0;
  assign out[463] = (in == 9'd463) ? 1'b1 : 1'b0;
  assign out[464] = (in == 9'd464) ? 1'b1 : 1'b0;
  assign out[465] = (in == 9'd465) ? 1'b1 : 1'b0;
  assign out[466] = (in == 9'd466) ? 1'b1 : 1'b0;
  assign out[467] = (in == 9'd467) ? 1'b1 : 1'b0;
  assign out[468] = (in == 9'd468) ? 1'b1 : 1'b0;
  assign out[469] = (in == 9'd469) ? 1'b1 : 1'b0;
  assign out[470] = (in == 9'd470) ? 1'b1 : 1'b0;
  assign out[471] = (in == 9'd471) ? 1'b1 : 1'b0;
  assign out[472] = (in == 9'd472) ? 1'b1 : 1'b0;
  assign out[473] = (in == 9'd473) ? 1'b1 : 1'b0;
  assign out[474] = (in == 9'd474) ? 1'b1 : 1'b0;
  assign out[475] = (in == 9'd475) ? 1'b1 : 1'b0;
  assign out[476] = (in == 9'd476) ? 1'b1 : 1'b0;
  assign out[477] = (in == 9'd477) ? 1'b1 : 1'b0;
  assign out[478] = (in == 9'd478) ? 1'b1 : 1'b0;
  assign out[479] = (in == 9'd479) ? 1'b1 : 1'b0;
  assign out[480] = (in == 9'd480) ? 1'b1 : 1'b0;
  assign out[481] = (in == 9'd481) ? 1'b1 : 1'b0;
  assign out[482] = (in == 9'd482) ? 1'b1 : 1'b0;
  assign out[483] = (in == 9'd483) ? 1'b1 : 1'b0;
  assign out[484] = (in == 9'd484) ? 1'b1 : 1'b0;
  assign out[485] = (in == 9'd485) ? 1'b1 : 1'b0;
  assign out[486] = (in == 9'd486) ? 1'b1 : 1'b0;
  assign out[487] = (in == 9'd487) ? 1'b1 : 1'b0;
  assign out[488] = (in == 9'd488) ? 1'b1 : 1'b0;
  assign out[489] = (in == 9'd489) ? 1'b1 : 1'b0;
  assign out[490] = (in == 9'd490) ? 1'b1 : 1'b0;
  assign out[491] = (in == 9'd491) ? 1'b1 : 1'b0;
  assign out[492] = (in == 9'd492) ? 1'b1 : 1'b0;
  assign out[493] = (in == 9'd493) ? 1'b1 : 1'b0;
  assign out[494] = (in == 9'd494) ? 1'b1 : 1'b0;
  assign out[495] = (in == 9'd495) ? 1'b1 : 1'b0;
  assign out[496] = (in == 9'd496) ? 1'b1 : 1'b0;
  assign out[497] = (in == 9'd497) ? 1'b1 : 1'b0;
  assign out[498] = (in == 9'd498) ? 1'b1 : 1'b0;
  assign out[499] = (in == 9'd499) ? 1'b1 : 1'b0;
  assign out[500] = (in == 9'd500) ? 1'b1 : 1'b0;
  assign out[501] = (in == 9'd501) ? 1'b1 : 1'b0;
  assign out[502] = (in == 9'd502) ? 1'b1 : 1'b0;
  assign out[503] = (in == 9'd503) ? 1'b1 : 1'b0;
  assign out[504] = (in == 9'd504) ? 1'b1 : 1'b0;
  assign out[505] = (in == 9'd505) ? 1'b1 : 1'b0;
  assign out[506] = (in == 9'd506) ? 1'b1 : 1'b0;
  assign out[507] = (in == 9'd507) ? 1'b1 : 1'b0;
  assign out[508] = (in == 9'd508) ? 1'b1 : 1'b0;
  assign out[509] = (in == 9'd509) ? 1'b1 : 1'b0;
  assign out[510] = (in == 9'd510) ? 1'b1 : 1'b0;
  assign out[511] = (in == 9'd511) ? 1'b1 : 1'b0;
endmodule
